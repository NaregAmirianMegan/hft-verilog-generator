`timescale 1ns / 1ps
`include "../fp_gt.v"

module fp_gt_tb();
    reg [31:0] F1;
    reg [31:0] F2;

    wire RESULT;

    fp_gt uut (.out(RESULT), .f1(F1), .f2(F2));

    initial begin
        $monitor("F1=%d, F2=%d, RESULT=%b", F1[30:0], F2[30:0], RESULT);
        $dumpfile("fp_gt.vcd");
        $dumpvars(0, fp_gt_tb);
        
        // Expect: 1
        F1 = 32'b01000001010000000000000000000000; // 12 
        F2 = 32'b11000001010000000000000000000000; // -12
        #100000;

        // Expect: 0
        F1 = 32'b11000001010000000000000000000000; // -12
        F2 = 32'b01000001010000000000000000000000; // 12
        #100000;

        // Expect: 0
        F1 = 32'b00000000000000000000000000000000; // 0
        F2 = 32'b01000001010101100110011001100110; // 13.4
        #100000;

        // Expect: 1
        F1 = 32'b01000001010101100110011001100110; // 13.4
        F2 = 32'b00000000000000000000000000000000; // 0
        #100000;

        // Expect: 1
        F1 = 32'b00000000000000000000000000000000; // 0
        F2 = 32'b11000001001000111010111000010100; // -10.23
        #100000;

        // Expect: 0
        F1 = 32'b11000001001000111010111000010100; // -10.23
        F2 = 32'b00000000000000000000000000000000; // 0
        #100000;

        // Expect: 1
        F1 = 32'b01000001110001000111101011100001; // 24.56
        F2 = 32'b01000001001000111010111000010100; // 10.23
        #100000;

        // Expect: 0
        F1 = 32'b01000001001000111010111000010100; // 10.23
        F2 = 32'b01000001110001000111101011100001; // 24.56
        #100000;

        // Expect: 0
        F1 = 32'b11000010000010100011110101110001; // -34.56
        F2 = 32'b11000001011001010111000010100100; // -14.34
        #100000;

        // Expect: 1
        F1 = 32'b11000001011001010111000010100100; // -14.34 
        F2 = 32'b11000010000010100011110101110001; // -34.56
        #100000;
        $finish;
    end

endmodule