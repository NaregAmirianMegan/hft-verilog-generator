// Using IEEE-754 Single Precision Float

module fp_gt (output out, input [31:0] f1, input [31:0] f2);

    reg out = 1'b0;

    always @ (*)
    begin 

    end
endmodule