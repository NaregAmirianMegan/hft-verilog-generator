`include "fp_gt.v"

module test(output out1, output out2, input [31:0] RSI);
  reg out1 = 1'b1;
  reg out2 = 1'b0;
